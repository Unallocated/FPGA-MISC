LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
 
ENTITY serial_tx_fifo_tb IS
END serial_tx_fifo_tb;
 
ARCHITECTURE behavior OF serial_tx_fifo_tb IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT serial_tx_fifo
    PORT(
         clk : IN  std_logic;
         rst : IN  std_logic;
         tx : OUT  std_logic;
         din : IN  std_logic_vector(7 downto 0);
         wr_clk : IN  std_logic;
         wr_en : IN  std_logic;
         full : OUT  std_logic;
         empty : OUT  std_logic
        );
    END COMPONENT;
    

   --Inputs
   signal clk : std_logic := '0';
   signal rst : std_logic := '0';
   signal din : std_logic_vector(7 downto 0) := (others => '0');
   signal wr_en : std_logic := '0';

 	--Outputs
   signal tx : std_logic;
   signal full : std_logic;
   signal empty : std_logic;

   -- Clock period definitions
   constant clk_period : time := 10 ns;
 

	 procedure send_data ( 
		data : std_logic_vector(7 downto 0);
		signal wr_en : out std_logic;
		signal din : out std_logic_vector(7 downto 0)) is
	 begin
		din <= data;
		wait for clk_period;
		wr_en <= '1';
		wait for clk_period;
		wr_en <= '0';
	 end send_data;

BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: serial_tx_fifo PORT MAP (
          clk => clk,
          rst => rst,
          tx => tx,
          din => din,
          wr_clk => clk,
          wr_en => wr_en,
          full => full,
          empty => empty
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 
   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	

      wait for clk_period*10;

			send_data(x"55", wr_en, din);
			send_data(x"FF", wr_en, din);
			send_data(x"7e", wr_en, din);
			send_data(x"28", wr_en, din);
			send_data(x"99", wr_en, din);
      -- insert stimulus here 

      wait;
   end process;

END;
