library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity eth3 is
end eth3;

architecture Behavioral of eth3 is

begin


end Behavioral;

