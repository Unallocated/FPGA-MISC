----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    18:18:23 12/06/2013 
-- Design Name: 
-- Module Name:    test2 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity test2 is
    Port ( clk : in  STD_LOGIC;
           rst : in  STD_LOGIC;
           sck : out  STD_LOGIC;
           so : out  STD_LOGIC;
           si : in  STD_LOGIC;
           cs : out  STD_LOGIC);
end test2;

architecture Behavioral of test2 is

begin


end Behavioral;

