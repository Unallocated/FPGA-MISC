library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity ram_test is
	Port(clk      : in    STD_LOGIC;
		 rst      : in    STD_LOGIC;
		 leds     : out   STD_LOGIC_VECTOR(7 downto 0);
		 ram_addr : out   STD_LOGIC_VECTOR(21 downto 0);
		 ram_data : inout STD_LOGIC_VECTOR(15 downto 0);
		 ram_clk  : out   STD_LOGIC;
--		 ram_wait : in    STD_LOGIC;
		 ram_lb   : out   STD_LOGIC;
		 ram_ub   : out   STD_LOGIC;
		 ram_ce   : out   STD_LOGIC;
		 ram_adv  : out   STD_LOGIC;
		 ram_cre  : out   STD_LOGIC;
		 ram_we   : out   STD_LOGIC;
		 ram_oe   : out   STD_LOGIC);
end ram_test;

architecture Behavioral of ram_test is
	COMPONENT clock_divider
		GENERIC(divide_by : integer);
		PORT(
			clk      : IN  std_logic;
			rst      : IN  std_logic;
			slow_clk : OUT std_logic
		);
	END COMPONENT;

	signal ram_state : integer   := 0;
	signal slow_clk  : std_logic := '0';
	
	type data_lut_t is array(0 to 255) of std_logic_vector(7 downto 0);
	constant data_lut : data_lut_t := ("10010011", "01011101", "11011111", "00101001", "00100100", "00000110", "00000010", "01100111", "01100010", "10111110", "00011000", "10111010", "11110110", "10010111", "11010100", "00110001", "01111010", "00011111", "00010011", "01100100", "01101001", "01000000", "01001101", "00010001", "00010101", "11011001", "10100101", "10010001", "01000110", "00110101", "00011111", "10001010", "01110000", "01001101", "01000011", "01100000", "01111011", "00110100", "10101010", "10111110", "01000001", "00101011", "01010000", "01101101", "10000001", "01001010", "01101010", "01101110", "10110101", "01100111", "10110010", "01001100", "01100001", "11101101", "11111100", "00110000", "00101110", "10111110", "01010110", "10010011", "10011101", "00011001", "00111100", "11110110", "10111011", "01111001", "00011101", "00111010", "01100010", "01101110", "11000011", "10111011", "11111001", "00110110", "00000111", "00010100", "00110011", "01011100", "00100111", "00100111", "10010100", "10110001", "00100110", "00101110", "01110101", "00101100", "01100110", "11011100", "00011010", "00101101", "11010011", "11110110", "11010010", "01001010", "01101111", "00010110", "01011111", "11100000", "10110100", "00001110", "01001001", "10111001", "11110101", "00101011", "10110110", "00011001", "00010000", "11100101", "01001101", "10001100", "10011110", "10100100", "11001101", "00000001", "10101011", "01001010", "11110101", "01010001", "00101011", "10001101", "10111101", "11010101", "10000010", "01010011", "10010100", "00011001", "01101001", "10110110", "01000011", "00110101", "10100011", "01000100", "10000001", "00110001", "10011101", "11001110", "10101100", "10000001", "00010011", "00111110", "00001011", "11101111", "10001010", "00111111", "00100000", "11101000", "10110011", "11010010", "11000101", "00011011", "01111110", "11111010", "01100110", "01011100", "00110100", "00001010", "01100011", "00100111", "01111111", "10010011", "01000001", "11111001", "01101011", "01100000", "01011110", "01010010", "01011011", "00011110", "10100000", "10111111", "11010000", "00101000", "01101011", "11010111", "01000010", "11001100", "11001110", "00001111", "10000001", "10001011", "10110111", "11100111", "10101101", "01000100", "10110001", "01110111", "11011110", "01101011", "01011111", "10111111", "01101101", "00110101", "11010001", "10001110", "11011001", "01001000", "01100001", "01000011", "00111000", "11101001", "11010000", "11111011", "11100001", "01010001", "10100101", "11000001", "01101011", "00001011", "00101110", "11010100", "11101010", "11100001", "00110110", "00100010", "10000100", "00100111", "00010110", "01011100", "11111011", "10010110", "00001011", "10000101", "10010100", "00000111", "00001001", "10011000", "10110000", "01011101", "00000101", "10001010", "11101011", "01010001", "11000000", "11101000", "01011000", "11100101", "11011101", "11100010", "01101000", "10000011", "10100111", "10100001", "10010111", "00100000", "11000111", "01100010", "00010100", "11010110", "10010111", "11011001", "00010001", "01110101", "10001000", "11101110", "00111100", "00100101");

begin

	ram_cre <= '0';

	process(slow_clk, rst)
		variable data : integer range 0 to (2**16) - 1 := 0;
	begin
		if (rst = '1') then
			data := 127;
			ram_state <= 0;
			leds <= (others => '0');
		elsif (rising_edge(slow_clk)) then
			case ram_state is
				when 0 =>
					ram_we <= '1';
					ram_adv <= '0';
					ram_clk <= '0';
					ram_oe <= '1';
					ram_addr <= "00" & x"0000f";
--					ram_data <= std_logic_vector(to_unsigned(data,16));
					ram_data <= data_lut(data) & data_lut(data);
				when 1 =>
					ram_ce <= '0';
				when 2 =>
					ram_lb <= '0';
					ram_ub <= '0';
				when 3 =>
					ram_we <= '0';
				when 4 =>
					ram_we <= '1';
				when 5 =>
					ram_data <= (others => '1');
				when 6 =>
					ram_data <= (others => 'Z');
				when 7 =>
					ram_ce <= '0';
					ram_oe <= '0';
				when 8 =>
					leds <= ram_data(7 downto 0);
					data := data + 1;
				when 9 =>
					ram_lb <= '1';
					ram_ub <= '1';
					ram_oe <= '1';
					ram_ce <= '1';
				when others =>
					null;
			end case;
			
			if(ram_state < 9) then
				ram_state <= ram_state + 1;
			else
				--null;
				ram_state <= 0;
			end if;
		end if;
	end process;

	clock_div : clock_divider
		Generic Map(divide_by => 1000000)
		PORT MAP(
			clk      => clk,
			rst      => rst,
			slow_clk => slow_clk
		);

end Behavioral;

